module top_tb;
    logic clk;

endmodule
module top ();

endmodule
